`timescale 1ns/1ps
module CLA_64bit(a,b,cin,sum,cout);
    input [63:0] a,b;
    input cin;
    output [63:0] sum;
    output cout;
    
    //---Write down your design here---//

    //---------------------------------//

endmodule
